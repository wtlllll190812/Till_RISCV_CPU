module Control (inst,aluSel);

endmodule 