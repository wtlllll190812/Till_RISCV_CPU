module cpu_top(inst,clk);
input reg[31:0] cpu_top;
// Control Control_inst()
endmodule